package apb_pkg;		
	import uvm_pkg::*;
	`include "uvm_macros.svh"
	`define no_of_transfer 2147483647
	`include "apb_defines.sv"
  	`include"apb_seq_items.sv"
	`include"apb_wseqs.sv"
	`include"apb_rseqs.sv"
	`include"apb_sequencer.sv"
	`include"apb_driver.sv"
	`include"apb_monitor.sv"
	`include"apb_agent.sv"
  	`include"apb_coverage.sv"
	`include"apb_scoreboard.sv"
	`include"apb_env.sv"
	`include"apb_base_test.sv"
endpackage