parameter ADDR_WIDTH = 32 ;
parameter DATA_WIDTH = 32;